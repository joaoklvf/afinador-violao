library verilog;
use verilog.vl_types.all;
entity afinador_violao_vlg_vec_tst is
end afinador_violao_vlg_vec_tst;
