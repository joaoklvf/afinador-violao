library verilog;
use verilog.vl_types.all;
entity oscilador_vlg_vec_tst is
end oscilador_vlg_vec_tst;
