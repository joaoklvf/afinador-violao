// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Fri May 24 21:51:00 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module UC (
    reset,clock,start);

    input reset;
    input clock;
    input start;
    tri0 reset;
    tri0 start;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter state1=0,state2=1,state3=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or start)
    begin
        if (reset) begin
            reg_fstate <= state1;
        end
        else begin
            case (fstate)
                state1: begin
                    if ((start == 1'b0))
                        reg_fstate <= state1;
                    else if ((start == 1'b1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    reg_fstate <= state3;
                end
                state3: begin
                    if ((start == 1'b1))
                        reg_fstate <= state3;
                    else if ((start == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;
                end
                default: begin
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // UC
